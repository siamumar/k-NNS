`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:56:45 09/23/2016
// Design Name:   k_nns_seq
// Module Name:   C:/Users/Rice/Dropbox/SFE/VerilogCodes/k_NNS/k_nns_seq_tb.v
// Project Name:  k_NNS
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: k_nns_seq
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module k_nns_seq_tb;

	parameter W = 32, K = 8;

	// Inputs
	reg clk;
	reg rst;
	wire [2*W-1:0] g_input;
	wire [2*W-1:0] e_init;

	// Outputs
	wire [2*W*K-1:0] o;

	// Instantiate the Unit Under Test (UUT)
	k_nns_seq #(.W(W), .K(K)) uut (
		.clk(clk), 
		.rst(rst), 
		.g_input(g_input), 
		.e_init(e_init), 
		.o(o)
	);
	
	reg [W-1:0] x1, y1, x2, y2;
	
	assign e_init[2*W-1:W]	=  x1;
	assign e_init[W-1:0]	=  y1;
	assign g_input[2*W-1:W]	=  x2;
	assign g_input[W-1:0]	=  y2;	
		
	wire signed [W-1:0] xR[K-1:0];	
	wire signed [W-1:0] yR[K-1:0];
	
	genvar i;
	
	generate
	for (i = K-1; i >= 0; i = i-1)
	begin:R_ASN
		assign xR[i] = o[W*(2*i+2)-1:W*(2*i+1)];
		assign yR[i] = o[W*(2*i+1)-1:W*2*i];
	end
	endgenerate
	
	integer j;

	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 1;
		x1 = 7305964; 
		y1 = 647733192; 
		x2 = 0;
		y2 = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		rst = 0;
		
		x1 = 0; 
		y1 = 0; 
		x2 = 1271116984; 
		y2 = 592265768; 
		#100; 
		x2 = -1145150946; 
		y2 = -2078249626; 
		#100; 
		x2 = 433099943; 
		y2 = 1700612176; 
		#100; 
		x2 = -1664461410; 
		y2 = 66035367; 
		#100; 
		x2 = 67712965; 
		y2 = 191220269; 
		#100; 
		x2 = 1451014718; 
		y2 = 457165803; 
		#100; 
		x2 = 1807279752; 
		y2 = 1118565038; 
		#100; 
		x2 = -7610985; 
		y2 = 1526203193; 
		#100; 
		x2 = -955152957; 
		y2 = -503076184; 
		#100; 
		x2 = 655068243; 
		y2 = -1783918151; 
		#100; 
		x2 = 1792284715; 
		y2 = 1004478169; 
		#100; 
		x2 = 42260131; 
		y2 = -721600322; 
		#100; 
		x2 = 2036636914; 
		y2 = 1459213141; 
		#100; 
		x2 = -1300177043; 
		y2 = -550944197; 
		#100; 
		x2 = -1669947778; 
		y2 = 1409673851; 
		#100; 
		x2 = -870356682; 
		y2 = -1389341909; 
		#100; 
		x2 = -444879002; 
		y2 = -1591200080; 
		#100; 
		x2 = -340351748; 
		y2 = 1631587562; 
		#100; 
		x2 = -809707173; 
		y2 = -1958165232; 
		#100; 
		x2 = 832550080; 
		y2 = 801956373; 
		#100; 
		x2 = -1752897128; 
		y2 = 1004046981; 
		#100; 
		x2 = -420526179; 
		y2 = -269842327; 
		#100; 
		x2 = -879691748; 
		y2 = -516087922; 
		#100; 
		x2 = -831090006; 
		y2 = 2060113017; 
		#100; 
		x2 = -1694102043; 
		y2 = -433819946; 
		#100; 
		x2 = 402986493; 
		y2 = -256895247; 
		#100; 
		x2 = -933178212; 
		y2 = -1473998899; 
		#100; 
		x2 = -1480811862; 
		y2 = -747177060; 
		#100; 
		x2 = -2144654692; 
		y2 = -798597935; 
		#100; 
		x2 = -929450606; 
		y2 = 1694367449; 
		#100; 
		x2 = 218231046; 
		y2 = -1086522876; 
		#100; 
		x2 = 1593012782; 
		y2 = -813127435; 
		#100; 
		x2 = -1966006568; 
		y2 = -391405060; 
		#100; 
		x2 = 1738267674; 
		y2 = 893399987; 
		#100; 
		x2 = -1584954230; 
		y2 = -1530564874; 
		#100; 
		x2 = 1433354918; 
		y2 = 1594816132; 
		#100; 
		x2 = 1290501843; 
		y2 = -1790331791; 
		#100; 
		x2 = 1794781328; 
		y2 = -164334733; 
		#100; 
		x2 = -1557768925; 
		y2 = -2016963785; 
		#100; 
		x2 = 20325149; 
		y2 = 1087488007; 
		#100; 
		x2 = -408200220; 
		y2 = 859176723; 
		#100; 
		x2 = -1401996890; 
		y2 = -1226160566; 
		#100; 
		x2 = 322911157; 
		y2 = 772684741; 
		#100; 
		x2 = 456202547; 
		y2 = 246070190; 
		#100; 
		x2 = -1226446206; 
		y2 = 1506154418; 
		#100; 
		x2 = 85608384; 
		y2 = 251536872; 
		#100; 
		x2 = 2101037054; 
		y2 = 1725604747; 
		#100; 
		x2 = -43314048; 
		y2 = -345668829; 
		#100; 
		x2 = 836974069; 
		y2 = -609334085; 
		#100; 
		x2 = -380440354; 
		y2 = -47298253; 
		#100; 
		x2 = -1998118686; 
		y2 = -1048134623; 
		#100; 
		x2 = -889781692; 
		y2 = 1843267974; 
		#100; 
		x2 = 1294682405; 
		y2 = -142778396; 
		#100; 
		x2 = -659268930; 
		y2 = -1056528237; 
		#100; 
		x2 = -1789644389; 
		y2 = -295414519; 
		#100; 
		x2 = 47701500; 
		y2 = 869859775; 
		#100; 
		x2 = -571946158; 
		y2 = -419490023; 
		#100; 
		x2 = 1028556641; 
		y2 = -1366486457; 
		#100; 
		x2 = 106258195; 
		y2 = 1530086893; 
		#100; 
		x2 = 1307907209; 
		y2 = 361641506; 
		#100; 
		x2 = 1361123149; 
		y2 = -542974994; 
		#100; 
		x2 = -1333709830; 
		y2 = -1195312820; 
		#100; 
		x2 = -1616224296; 
		y2 = -1206911074; 
		#100; 
		x2 = 1378669379; 
		y2 = 95487616; 
		#100;
		
		for (j = 0; j < K; j = j+1)
			$display("%d\t%d", xR[j], yR[j]);
	end
	
always begin
	#50;
	clk = ~clk;
end


      
endmodule

